LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY sbox IS
PORT(
    sbox_in    :	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
    sbox_out   :	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END sbox;

ARCHITECTURE beh OF sbox IS
    
BEGIN
--s box table
WITH sbox_in(7 DOWNTO 0) SELECT
    
sbox_out(7 DOWNTO 0) <= 
		    --first row
		    "01100011" WHEN "00000000", --(X"63")
		    "01111100" WHEN "00000001", --(X"7C") 
		    "01110111" WHEN "00000010", --(X"77")
		    "01111011" WHEN "00000011", --(X"7B")
		    "11110010" WHEN "00000100", --(X"F2")
		    "01101011" WHEN "00000101", --(X"6B")
		    "01101111" WHEN "00000110", --(X"6F") 
		    "11000101" WHEN "00000111", --(X"C5") 
		    "00110000" WHEN "00001000", --(X"30") 
		    "00000001" WHEN "00001001", --(X"01") 
		    "01100111" WHEN "00001010", --(X"67") 
		    "00101011" WHEN "00001011", --(X"2B") 
		    "11111110" WHEN "00001100", --(X"FE") 
		    "11010111" WHEN "00001101", --(X"D7") 
		    "10101011" WHEN "00001110", --(X"AB") 
		    "01110110" WHEN "00001111", --(X"76") 
		    --second row
		    "11001010" WHEN "00010000", --(X"CA") 
		    "10000010" WHEN "00010001", --(X"82")
		    "11001001" WHEN "00010010", --(X"C9")
		    "01111101" WHEN "00010011", --(X"7D")
		    "11111010" WHEN "00010100", --(X"FA")
		    "01011001" WHEN "00010101", --(X"59")
		    "01000111" WHEN "00010110", --(X"47")
		    "11110000" WHEN "00010111", --(X"F0")
		    "10101101" WHEN "00011000", --(X"AD")
		    "11010100" WHEN "00011001", --(X"D4")
		    "10100010" WHEN "00011010", --(X"A2")
		    "10101111" WHEN "00011011", --(X"AF")
		    "10011100" WHEN "00011100", --(X"9C")
		    "10100100" WHEN "00011101", --(X"A4")
		    "01110010" WHEN "00011110", --(X"72")
		    "11000000" WHEN "00011111", --(X"C0")
		    --third row
		    "10110111" WHEN "00100000", --(X"B7")
		    "11111101" WHEN "00100001", --(X"FD")
		    "10010011" WHEN "00100010", --(X"93")
		    "00100110" WHEN "00100011", --(X"26")
		    "00110110" WHEN "00100100", --(X"36")
		    "00111111" WHEN "00100101", --(X"3F")
		    "11110111" WHEN "00100110", --(X"F7")
		    "11001100" WHEN "00100111", --(X"CC")
		    "00110100" WHEN "00101000", --(X"34")
		    "10100101" WHEN "00101001", --(X"A5")
		    "11100101" WHEN "00101010", --(X"E5")
		    "11110001" WHEN "00101011", --(X"F1")
		    "01110001" WHEN "00101100", --(X"71")
		    "11011000" WHEN "00101101", --(X"D8")
		    "00110001" WHEN "00101110", --(X"31")
		    "00010101" WHEN "00101111", --(X"15")
		    --forth row
		    "00000100" WHEN "00110000", --(X"04")
		    "11000111" WHEN "00110001", --(X"C7")
		    "00100011" WHEN "00110010", --(X"23")
		    "11000011" WHEN "00110011", --(X"C3")
		    "00011000" WHEN "00110100", --(X"18")
		    "10010110" WHEN "00110101", --(X"96")
		    "00000101" WHEN "00110110", --(X"05")
		    "10011010" WHEN "00110111", --(X"9A")
		    "00000111" WHEN "00111000", --(X"07")
		    "00010010" WHEN "00111001", --(X"12")
		    "10000000" WHEN "00111010", --(X"80")
		    "11100010" WHEN "00111011", --(X"E2")
		    "11101011" WHEN "00111100", --(X"EB")
		    "00100111" WHEN "00111101", --(X"27")
		    "10110010" WHEN "00111110", --(X"B2")
		    "01110101" WHEN "00111111", --(X"75")
		    --fifth row
		    "00001001" WHEN "01000000", --(X"09") 
		    "10000011" WHEN "01000001", --(X"83") 
		    "00101100" WHEN "01000010", --(X"2C") 
		    "00011010" WHEN "01000011", --(X"1A") 
		    "00011011" WHEN "01000100", --(X"1B") 
		    "01101110" WHEN "01000101", --(X"6E") 
		    "01011010" WHEN "01000110", --(X"5A") 
		    "10100000" WHEN "01000111", --(X"A0") 
		    "01010010" WHEN "01001000", --(X"52") 
		    "00111011" WHEN "01001001", --(X"3B") 
		    "11010110" WHEN "01001010", --(X"D6") 
		    "10110011" WHEN "01001011", --(X"B3") 
		    "00101001" WHEN "01001100", --(X"29") 
		    "11100011" WHEN "01001101", --(X"E3") 
		    "00101111" WHEN "01001110", --(X"2F") 
		    "10000100" WHEN "01001111", --(X"84") 
		    --sixth row
		    "01010011" WHEN "01010000", --(X"53") 
		    "11010001" WHEN "01010001", --(X"D1") 
		    "00000000" WHEN "01010010", --(X"00") 
		    "11101101" WHEN "01010011", --(X"ED") 
		    "00100000" WHEN "01010100", --(X"20") 
		    "11111100" WHEN "01010101", --(X"FC") 
		    "10110001" WHEN "01010110", --(X"B1") 
		    "01011011" WHEN "01010111", --(X"5B") 
		    "01101010" WHEN "01011000", --(X"6A") 
		    "11001011" WHEN "01011001", --(X"CB") 
		    "10111110" WHEN "01011010", --(X"BE") 
		    "00111001" WHEN "01011011", --(X"39") 
		    "01001010" WHEN "01011100", --(X"4A") 
		    "01001100" WHEN "01011101", --(X"4C") 
		    "01011000" WHEN "01011110", --(X"58")
		    "11001111" WHEN "01011111", --(X"CF") 
		    --seventh row
		    "11010000" WHEN "01100000", --(X"D0") 
		    "11101111" WHEN "01100001", --(X"EF") 
		    "10101010" WHEN "01100010", --(X"AA") 
		    "11111011" WHEN "01100011", --(X"FB") 
		    "01000011" WHEN "01100100", --(X"43") 
		    "01001101" WHEN "01100101", --(X"4D") 
		    "00110011" WHEN "01100110", --(X"33") 
		    "10000101" WHEN "01100111", --(X"85") 
		    "01000101" WHEN "01101000", --(X"45") 
		    "11111001" WHEN "01101001", --(X"F9") 
		    "00000010" WHEN "01101010", --(X"02") 
		    "01111111" WHEN "01101011", --(X"7F") 
		    "01010000" WHEN "01101100", --(X"50") 
		    "00111100" WHEN "01101101", --(X"3C") 
		    "10011111" WHEN "01101110", --(X"9F") 
		    "10101000" WHEN "01101111", --(X"A8") 
		    --eighth row
		    "01010001" WHEN "01110000", --(X"51")
		    "10100011" WHEN "01110001", --(X"A3")
		    "01000000" WHEN "01110010", --(X"40")
		    "10001111" WHEN "01110011", --(X"8F")
		    "10010010" WHEN "01110100", --(X"92")
		    "10011101" WHEN "01110101", --(X"9D")
		    "00111000" WHEN "01110110", --(X"38")
		    "11110101" WHEN "01110111", --(X"F5")
		    "10111100" WHEN "01111000", --(X"BC")
		    "10110110" WHEN "01111001", --(X"B6")
		    "11011010" WHEN "01111010", --(X"DA")
		    "00100001" WHEN "01111011", --(X"21")
		    "00010000" WHEN "01111100", --(X"10")
		    "11111111" WHEN "01111101", --(X"FF")
		    "11110011" WHEN "01111110", --(X"F3")
		    "11010010" WHEN "01111111", --(X"D2")
		    --ninth row
		    "11001101" WHEN "10000000", --(X"CD") 
		    "00001100" WHEN "10000001", --(X"0C") 
		    "00010011" WHEN "10000010", --(X"13") 
		    "11101100" WHEN "10000011", --(X"EC") 
		    "01011111" WHEN "10000100", --(X"5F") 
		    "10010111" WHEN "10000101", --(X"97") 
		    "01000100" WHEN "10000110", --(X"44") 
		    "00010111" WHEN "10000111", --(X"17") 
		    "11000100" WHEN "10001000", --(X"C4") 
		    "10100111" WHEN "10001001", --(X"A7") 
		    "01111110" WHEN "10001010", --(X"7E") 
		    "00111101" WHEN "10001011", --(X"3D") 
		    "01100100" WHEN "10001100", --(X"64") 
		    "01011101" WHEN "10001101", --(X"5D") 
		    "00011001" WHEN "10001110", --(X"19") 
		    "01110011" WHEN "10001111", --(X"73") 
		    --tenth row
		    "01100000" WHEN "10010000", --(X"60") 
		    "10000001" WHEN "10010001", --(X"81") 
		    "01001111" WHEN "10010010", --(X"4F") 
		    "11011100" WHEN "10010011", --(X"DC") 
		    "00100010" WHEN "10010100", --(X"22") 
		    "00101010" WHEN "10010101", --(X"2A") 
		    "10010000" WHEN "10010110", --(X"90") 
		    "10001000" WHEN "10010111", --(X"88") 
		    "01000110" WHEN "10011000", --(X"46") 
		    "11101110" WHEN "10011001", --(X"EE") 
		    "10111000" WHEN "10011010", --(X"B8")
		    "00010100" WHEN "10011011", --(X"14") 
		    "11011110" WHEN "10011100", --(X"DE")
		    "01011110" WHEN "10011101", --(X"5E") 
		    "00001011" WHEN "10011110", --(X"0B")
		    "11011011" WHEN "10011111", --(X"DB") 
		    --eleventh row
		    "11100000" WHEN "10100000", --(X"E0") 
		    "00110010" WHEN "10100001", --(X"32") 
		    "00111010" WHEN "10100010", --(X"3A") 
		    "00001010" WHEN "10100011", --(X"0A") 
		    "01001001" WHEN "10100100", --(X"49") 
		    "00000110" WHEN "10100101", --(X"06") 
		    "00100100" WHEN "10100110", --(X"24") 
		    "01011100" WHEN "10100111", --(X"5C") 
		    "11000010" WHEN "10101000", --(X"C2") 
		    "11010011" WHEN "10101001", --(X"D3") 
		    "10101100" WHEN "10101010", --(X"AC") 
		    "01100010" WHEN "10101011", --(X"62") 
		    "10010001" WHEN "10101100", --(X"91") 
		    "10010101" WHEN "10101101", --(X"95") 
		    "11100100" WHEN "10101110", --(X"E4") 
		    "01111001" WHEN "10101111", --(X"79") 
		    --twelveth row
		    "11100111" WHEN "10110000", --(X"E7") 
		    "11001000" WHEN "10110001", --(X"C8") 
		    "00110111" WHEN "10110010", --(X"37") 
		    "01101101" WHEN "10110011", --(X"6D") 
		    "10001101" WHEN "10110100", --(X"8D") 
		    "11010101" WHEN "10110101", --(X"D5") 
		    "01001110" WHEN "10110110", --(X"4E") 
		    "10101001" WHEN "10110111", --(X"A9") 
		    "01101100" WHEN "10111000", --(X"6C") 
		    "01010110" WHEN "10111001", --(X"56") 
		    "11110100" WHEN "10111010", --(X"F4") 
		    "11101010" WHEN "10111011", --(X"EA") 
		    "01100101" WHEN "10111100", --(X"65") 
		    "01111010" WHEN "10111101", --(X"7A") 
		    "10101110" WHEN "10111110", --(X"AE") 
		    "00001000" WHEN "10111111", --(X"08") 
		    --thirteenth row
		    "10111010" WHEN "11000000", --(X"BA") 
		    "01111000" WHEN "11000001", --(X"78") 
		    "00100101" WHEN "11000010", --(X"25") 
		    "00101110" WHEN "11000011", --(X"2E") 
		    "00011100" WHEN "11000100", --(X"1C")
		    "10100110" WHEN "11000101", --(X"A6") 
		    "10110100" WHEN "11000110", --(X"B4") 
		    "11000110" WHEN "11000111", --(X"C6") 
		    "11101000" WHEN "11001000", --(X"E8") 
		    "11011101" WHEN "11001001", --(X"DD") 
		    "01110100" WHEN "11001010", --(X"74") 
		    "00011111" WHEN "11001011", --(X"1F") 
		    "01001011" WHEN "11001100", --(X"4B") 
		    "10111101" WHEN "11001101", --(X"BD") 
		    "10001011" WHEN "11001110", --(X"8B") 
		    "10001010" WHEN "11001111", --(X"8A") 
		    --forteenth row
		    "01110000" WHEN "11010000", --(X"70") 
		    "00111110" WHEN "11010001", --(X"3E") 
		    "10110101" WHEN "11010010", --(X"B5") 
		    "01100110" WHEN "11010011", --(X"66") 
		    "01001000" WHEN "11010100", --(X"48") 
		    "00000011" WHEN "11010101", --(X"03") 
		    "11110110" WHEN "11010110", --(X"F6") 
		    "00001110" WHEN "11010111", --(X"0E") 
		    "01100001" WHEN "11011000", --(X"61") 
		    "00110101" WHEN "11011001", --(X"35") 
		    "01010111" WHEN "11011010", --(X"57") 
		    "10111001" WHEN "11011011", --(X"B9") 
		    "10000110" WHEN "11011100", --(X"86") 
		    "11000001" WHEN "11011101", --(X"C1") 
		    "00011101" WHEN "11011110", --(X"1D") 
		    "10011110" WHEN "11011111", --(X"9E") 
		    --fifteenth row
		    "11100001" WHEN "11100000", --(X"E1") 
		    "11111000" WHEN "11100001", --(X"F8") 
		    "10011000" WHEN "11100010", --(X"98") 
		    "00010001" WHEN "11100011", --(X"11") 
		    "01101001" WHEN "11100100", --(X"69") 
		    "11011001" WHEN "11100101", --(X"D9") 
		    "10001110" WHEN "11100110", --(X"8E") 
		    "10010100" WHEN "11100111", --(X"94") 
		    "10011011" WHEN "11101000", --(X"9B") 
		    "00011110" WHEN "11101001", --(X"1E") 
		    "10000111" WHEN "11101010", --(X"87") 
		    "11101001" WHEN "11101011", --(X"E9") 
		    "11001110" WHEN "11101100", --(X"CE") 
		    "01010101" WHEN "11101101", --(X"55") 
		    "00101000" WHEN "11101110", --(X"28") 
		    "11011111" WHEN "11101111", --(X"DF") 
		    --sixteenth row
		    "10001100" WHEN "11110000", --(X"8C") 
		    "10100001" WHEN "11110001", --(X"A1") 
		    "10001001" WHEN "11110010", --(X"89") 
		    "00001101" WHEN "11110011", --(X"0D") 
		    "10111111" WHEN "11110100", --(X"BF") 
		    "11100110" WHEN "11110101", --(X"E6") 
		    "01000010" WHEN "11110110", --(X"42") 
		    "01101000" WHEN "11110111", --(X"68") 
		    "01000001" WHEN "11111000", --(X"41") 
		    "10011001" WHEN "11111001", --(X"99") 
		    "00101101" WHEN "11111010", --(X"2D") 
		    "00001111" WHEN "11111011", --(X"0F") 
		    "10110000" WHEN "11111100", --(X"B0") 
		    "01010100" WHEN "11111101", --(X"54") 
		    "10111011" WHEN "11111110", --(X"BB") 
		    "00010110" WHEN "11111111", --(X"16") 
		    
		    "XXXXXXXX" WHEN OTHERS;
END beh;			    
			    
